// megafunction wizard: %LPM_DIVIDE%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: LPM_DIVIDE 

// ============================================================
// File Name: div_int.v
// Megafunction Name(s):
// 			LPM_DIVIDE
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 17.1.0 Build 590 10/25/2017 SJ Lite Edition
// ************************************************************

//Copyright (C) 2017  Intel Corporation. All rights reserved.
//Your use of Intel Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Intel Program License 
//Subscription Agreement, the Intel Quartus Prime License Agreement,
//the Intel FPGA IP License Agreement, or other applicable license
//agreement, including, without limitation, that your use is for
//the sole purpose of programming logic devices manufactured by
//Intel and sold by Intel or its authorized distributors.  Please
//refer to the applicable agreement for further details.

module div_int (
	denom,
	numer,
	quotient,
	remain);

	input	[5:0]  denom;
	input	[5:0]  numer;
	output	[5:0]  quotient;
	output	[5:0]  remain;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: PRIVATE: PRIVATE_LPM_REMAINDERPOSITIVE STRING "TRUE"
// Retrieval info: PRIVATE: PRIVATE_MAXIMIZE_SPEED NUMERIC "6"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: USING_PIPELINE NUMERIC "0"
// Retrieval info: PRIVATE: VERSION_NUMBER NUMERIC "2"
// Retrieval info: PRIVATE: new_diagram STRING "1"
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: CONSTANT: LPM_DREPRESENTATION STRING "UNSIGNED"
// Retrieval info: CONSTANT: LPM_HINT STRING "MAXIMIZE_SPEED=6,LPM_REMAINDERPOSITIVE=TRUE"
// Retrieval info: CONSTANT: LPM_NREPRESENTATION STRING "UNSIGNED"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_DIVIDE"
// Retrieval info: CONSTANT: LPM_WIDTHD NUMERIC "6"
// Retrieval info: CONSTANT: LPM_WIDTHN NUMERIC "6"
// Retrieval info: USED_PORT: denom 0 0 6 0 INPUT NODEFVAL "denom[5..0]"
// Retrieval info: USED_PORT: numer 0 0 6 0 INPUT NODEFVAL "numer[5..0]"
// Retrieval info: USED_PORT: quotient 0 0 6 0 OUTPUT NODEFVAL "quotient[5..0]"
// Retrieval info: USED_PORT: remain 0 0 6 0 OUTPUT NODEFVAL "remain[5..0]"
// Retrieval info: CONNECT: @denom 0 0 6 0 denom 0 0 6 0
// Retrieval info: CONNECT: @numer 0 0 6 0 numer 0 0 6 0
// Retrieval info: CONNECT: quotient 0 0 6 0 @quotient 0 0 6 0
// Retrieval info: CONNECT: remain 0 0 6 0 @remain 0 0 6 0
// Retrieval info: GEN_FILE: TYPE_NORMAL div_int.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL div_int.inc TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL div_int.cmp TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL div_int.bsf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL div_int_inst.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL div_int_bb.v TRUE
// Retrieval info: LIB_FILE: lpm
