
module DE0_CV_golden_top (

);
endmodule 
